`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Bucknell University 
// Engineer: Yifan Ge, Alex Thompson
// 
// Create Date:    16:57:48 04/21/2012 
// Design Name: Memory Game font
// Module Name:    font_rom 
// Project Name: Project 3 ELEC 340
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module font_rom(
	 input wire clk,
	 input wire [8:0] addr,
	 output reg [23:0] data
    );
	 
	 // Registers used to access font ROM
	 reg [8:0] addr_reg;
	 reg [23:0] data_reg;
	 
	 always @ (posedge clk)
		addr_reg <= addr;
	 
	 // Font ROM
	 always @ *
		case (addr_reg)
			// Zero
			9'h000 : data = 24'b000011111111111111110000;
			9'h001 : data = 24'b000111111111111111111000;
			9'h002 : data = 24'b001111111111111111111100;
			9'h003 : data = 24'b011111111111111111111110;
			9'h004 : data = 24'b111111100000000001111111;
			9'h005 : data = 24'b111111000000000000111111;
			9'h006 : data = 24'b111110000000000000111111;
			9'h007 : data = 24'b111100000000000001111111;
			9'h008 : data = 24'b111100000000000011111111;
			9'h009 : data = 24'b111100000000000111111111;
			9'h00a : data = 24'b111100000000001111111111;
			9'h00b : data = 24'b111100000000011111111111;
			9'h00c : data = 24'b111100000000111111101111;
			9'h00d : data = 24'b111100000001111111001111;
			9'h00e : data = 24'b111100000011111110001111;
			9'h00f : data = 24'b111100000111111100001111;
			9'h010 : data = 24'b111100001111111000001111;
			9'h011 : data = 24'b111100011111110000001111;
			9'h012 : data = 24'b111100111111100000001111;
			9'h013 : data = 24'b111101111111000000001111;
			9'h014 : data = 24'b111111111110000000001111;
			9'h015 : data = 24'b111111111100000000001111;
			9'h016 : data = 24'b111111111000000000001111;
			9'h017 : data = 24'b111111110000000000001111;
			9'h018 : data = 24'b111111100000000000001111;
			9'h019 : data = 24'b111111000000000000011111;
			9'h01a : data = 24'b111111000000000000111111;
			9'h01b : data = 24'b111111100000000001111111;
			9'h01c : data = 24'b011111111111111111111110;
			9'h01d : data = 24'b001111111111111111111100;
			9'h01e : data = 24'b000111111111111111111000;
			9'h01f : data = 24'b000011111111111111110000;
			
			// One
			9'h020 : data = 24'b000000000000111100000000;
			9'h021 : data = 24'b000000000001111100000000;
			9'h022 : data = 24'b000000000011111100000000;
			9'h023 : data = 24'b000000000111111100000000;
			9'h024 : data = 24'b000000001111111100000000;
			9'h025 : data = 24'b000000011111111100000000;
			9'h026 : data = 24'b000000111110111100000000;
			9'h027 : data = 24'b000001111100111100000000;
			9'h028 : data = 24'b000011111000111100000000;
			9'h029 : data = 24'b000011110000111100000000;
			9'h02a : data = 24'b000011100000111100000000;
			9'h02b : data = 24'b000011000000111100000000;
			9'h02c : data = 24'b000000000000111100000000;
			9'h02d : data = 24'b000000000000111100000000;
			9'h02e : data = 24'b000000000000111100000000;
			9'h02f : data = 24'b000000000000111100000000;
			9'h030 : data = 24'b000000000000111100000000;
			9'h031 : data = 24'b000000000000111100000000;
			9'h032 : data = 24'b000000000000111100000000;
			9'h033 : data = 24'b000000000000111100000000;
			9'h034 : data = 24'b000000000000111100000000;
			9'h035 : data = 24'b000000000000111100000000;
			9'h036 : data = 24'b000000000000111100000000;
			9'h037 : data = 24'b000000000000111100000000;
			9'h038 : data = 24'b000000000000111100000000;
			9'h039 : data = 24'b000000000000111100000000;
			9'h03a : data = 24'b000000000000111100000000;
			9'h03b : data = 24'b000000000000111100000000;
			9'h03c : data = 24'b000011111111111111111111;
			9'h03d : data = 24'b000011111111111111111111;
			9'h03e : data = 24'b000011111111111111111111;
			9'h03f : data = 24'b000011111111111111111111;
			
			// Two
			9'h040 : data = 24'b000111111111111111110000;
			9'h041 : data = 24'b001111111111111111111000;
			9'h042 : data = 24'b011111111111111111111100;
			9'h043 : data = 24'b111111111111111111111110;
			9'h044 : data = 24'b111111100000000001111111;
			9'h045 : data = 24'b111111000000000000111111;
			9'h046 : data = 24'b111110000000000000011111;
			9'h047 : data = 24'b111110000000000000001111;
			9'h048 : data = 24'b000000000000000000001111;
			9'h049 : data = 24'b000000000000000000011111;
			9'h04a : data = 24'b000000000000000000111111;
			9'h04b : data = 24'b000000000000000001111111;
			9'h04c : data = 24'b000000000000000011111110;
			9'h04d : data = 24'b000000000000000111111100;
			9'h04e : data = 24'b000000000000001111111000;
			9'h04f : data = 24'b000000000000011111110000;
			9'h050 : data = 24'b000000000000111111100000;
			9'h051 : data = 24'b000000000001111111000000;
			9'h052 : data = 24'b000000000011111110000000;
			9'h053 : data = 24'b000000000111111100000000;
			9'h054 : data = 24'b000000001111111000000000;
			9'h055 : data = 24'b000000011111110000000000;
			9'h056 : data = 24'b000000111111100000000000;
			9'h057 : data = 24'b000001111111000000000000;
			9'h058 : data = 24'b000011111110000000000000;
			9'h059 : data = 24'b000111111100000000000000;
			9'h05a : data = 24'b001111111000000000000000;
			9'h05b : data = 24'b011111110000000000000000;
			9'h05c : data = 24'b111111111111111111111111;
			9'h05d : data = 24'b111111111111111111111111;
			9'h05e : data = 24'b111111111111111111111111;
			9'h05f : data = 24'b111111111111111111111111;
			
			// Three
			9'h060 : data = 24'b000111111111111111110000;
			9'h061 : data = 24'b001111111111111111111000;
			9'h062 : data = 24'b011111111111111111111100;
			9'h063 : data = 24'b111111111111111111111110;
			9'h064 : data = 24'b111111100000000001111111;
			9'h065 : data = 24'b111111000000000000111111;
			9'h066 : data = 24'b111110000000000000011111;
			9'h067 : data = 24'b111110000000000000001111;
			9'h068 : data = 24'b000000000000000000001111;
			9'h069 : data = 24'b000000000000000000001111;
			9'h06a : data = 24'b000000000000000000001111;
			9'h06b : data = 24'b000000000000000000011111;
			9'h06c : data = 24'b000000000000000000111111;
			9'h06d : data = 24'b000000000000000001111110;
			9'h06e : data = 24'b000011111111111111111100;
			9'h06f : data = 24'b000011111111111111111000;
			9'h070 : data = 24'b000011111111111111111100;
			9'h071 : data = 24'b000011111111111111111110;
			9'h072 : data = 24'b000000000000000001111111;
			9'h073 : data = 24'b000000000000000000111111;
			9'h074 : data = 24'b000000000000000000011111;
			9'h075 : data = 24'b000000000000000000001111;
			9'h076 : data = 24'b000000000000000000001111;
			9'h077 : data = 24'b000000000000000000001111;
			9'h078 : data = 24'b111110000000000000001111;
			9'h079 : data = 24'b111110000000000000011111;
			9'h07a : data = 24'b111111000000000000111111;
			9'h07b : data = 24'b111111100000000001111111;
			9'h07c : data = 24'b111111111111111111111110;
			9'h07d : data = 24'b011111111111111111111100;
			9'h07e : data = 24'b001111111111111111111000;
			9'h07f : data = 24'b000111111111111111110000;
			
			// Four
			9'h080 : data = 24'b000000000000000011110000;
			9'h081 : data = 24'b000000000000000111110000;
			9'h082 : data = 24'b000000000000001111110000;
			9'h083 : data = 24'b000000000000011111110000;
			9'h084 : data = 24'b000000000000111111110000;
			9'h085 : data = 24'b000000000001111111110000;
			9'h086 : data = 24'b000000000011111111110000;
			9'h087 : data = 24'b000000000111111111110000;
			9'h088 : data = 24'b000000001111111011110000;
			9'h089 : data = 24'b000000011111110011110000;
			9'h08a : data = 24'b000000111111100011110000;
			9'h08b : data = 24'b000001111111000011110000;
			9'h08c : data = 24'b000011111110000011110000;
			9'h08d : data = 24'b000111111100000011110000;
			9'h08e : data = 24'b001111111000000011110000;
			9'h08f : data = 24'b011111110000000011110000;
			9'h090 : data = 24'b111111111111111111111111;
			9'h091 : data = 24'b111111111111111111111111;
			9'h092 : data = 24'b111111111111111111111111;
			9'h093 : data = 24'b111111111111111111111111;
			9'h094 : data = 24'b000000000000000011110000;
			9'h095 : data = 24'b000000000000000011110000;
			9'h096 : data = 24'b000000000000000011110000;
			9'h097 : data = 24'b000000000000000011110000;
			9'h098 : data = 24'b000000000000000011110000;
			9'h099 : data = 24'b000000000000000011110000;
			9'h09a : data = 24'b000000000000000011110000;
			9'h09b : data = 24'b000000000000000011110000;
			9'h09c : data = 24'b000000000000111111111111;
			9'h09d : data = 24'b000000000000111111111111;
			9'h09e : data = 24'b000000000000111111111111;
			9'h09f : data = 24'b000000000000111111111111;
			
			// Five
			9'h0a0 : data = 24'b111111111111111111111111;
			9'h0a1 : data = 24'b111111111111111111111111;
			9'h0a2 : data = 24'b111111111111111111111111;
			9'h0a3 : data = 24'b111111111111111111111111;
			9'h0a4 : data = 24'b111100000000000000000000;
			9'h0a5 : data = 24'b111100000000000000000000;
			9'h0a6 : data = 24'b111100000000000000000000;
			9'h0a7 : data = 24'b111100000000000000000000;
			9'h0a8 : data = 24'b111100000000000000000000;
			9'h0a9 : data = 24'b111100000000000000000000;
			9'h0aa : data = 24'b111100000000000000000000;
			9'h0ab : data = 24'b111100000000000000000000;
			9'h0ac : data = 24'b111111111111111111111000;
			9'h0ad : data = 24'b111111111111111111111100;
			9'h0ae : data = 24'b111111111111111111111110;
			9'h0af : data = 24'b111111111111111111111111;
			9'h0b0 : data = 24'b000000000000000001111111;
			9'h0b1 : data = 24'b000000000000000000111111;
			9'h0b2 : data = 24'b000000000000000000011111;
			9'h0b3 : data = 24'b000000000000000000001111;
			9'h0b4 : data = 24'b000000000000000000001111;
			9'h0b5 : data = 24'b000000000000000000001111;
			9'h0b6 : data = 24'b000000000000000000001111;
			9'h0b7 : data = 24'b000000000000000000001111;
			9'h0b8 : data = 24'b111110000000000000001111;
			9'h0b9 : data = 24'b111110000000000000011111;
			9'h0ba : data = 24'b111111000000000000111111;
			9'h0bb : data = 24'b111111100000000001111111;
			9'h0bc : data = 24'b111111111111111111111111;
			9'h0bd : data = 24'b011111111111111111111110;
			9'h0be : data = 24'b001111111111111111111100;
			9'h0bf : data = 24'b000111111111111111111000;
			
			// Six
			9'h0c0 : data = 24'b000111111111111111111000;
			9'h0c1 : data = 24'b001111111111111111111100;
			9'h0c2 : data = 24'b011111111111111111111110;
			9'h0c3 : data = 24'b111111111111111111111111;
			9'h0c4 : data = 24'b111111100000000001111111;
			9'h0c5 : data = 24'b111111000000000000111111;
			9'h0c6 : data = 24'b111110000000000000011111;
			9'h0c7 : data = 24'b111100000000000000011111;
			9'h0c8 : data = 24'b111100000000000000000000;
			9'h0c9 : data = 24'b111100000000000000000000;
			9'h0ca : data = 24'b111100000000000000000000;
			9'h0cb : data = 24'b111100000000000000000000;
			9'h0cc : data = 24'b111111111111111111111000;
			9'h0cd : data = 24'b111111111111111111111100;
			9'h0ce : data = 24'b111111111111111111111110;
			9'h0cf : data = 24'b111111111111111111111111;
			9'h0d0 : data = 24'b111111100000000001111111;
			9'h0d1 : data = 24'b111111000000000000111111;
			9'h0d2 : data = 24'b111110000000000000011111;
			9'h0d3 : data = 24'b111100000000000000001111;
			9'h0d4 : data = 24'b111100000000000000001111;
			9'h0d5 : data = 24'b111100000000000000001111;
			9'h0d6 : data = 24'b111100000000000000001111;
			9'h0d7 : data = 24'b111100000000000000001111;
			9'h0d8 : data = 24'b111100000000000000001111;
			9'h0d9 : data = 24'b111110000000000000011111;
			9'h0da : data = 24'b111111000000000000111111;
			9'h0db : data = 24'b111111100000000001111111;
			9'h0dc : data = 24'b111111111111111111111111;
			9'h0dd : data = 24'b011111111111111111111110;
			9'h0de : data = 24'b001111111111111111111100;
			9'h0df : data = 24'b000111111111111111111000;
			
			// Seven
			9'h0e0 : data = 24'b111111111111111111111111;
			9'h0e1 : data = 24'b111111111111111111111111;
			9'h0e2 : data = 24'b111111111111111111111111;
			9'h0e3 : data = 24'b111111111111111111111111;
			9'h0e4 : data = 24'b000000000000000000001111;
			9'h0e5 : data = 24'b000000000000000000001111;
			9'h0e6 : data = 24'b000000000000000000001111;
			9'h0e7 : data = 24'b000000000000000000001111;
			9'h0e8 : data = 24'b000000000000000000001111;
			9'h0e9 : data = 24'b000000000000000000011111;
			9'h0ea : data = 24'b000000000000000000111111;
			9'h0eb : data = 24'b000000000000000001111111;
			9'h0ec : data = 24'b000000000000000011111110;
			9'h0ed : data = 24'b000000000000000111111100;
			9'h0ee : data = 24'b000000000000001111111000;
			9'h0ef : data = 24'b000000000000011111110000;
			9'h0f0 : data = 24'b000000000000111111100000;
			9'h0f1 : data = 24'b000000000001111111000000;
			9'h0f2 : data = 24'b000000000011111110000000;
			9'h0f3 : data = 24'b000000000111111100000000;
			9'h0f4 : data = 24'b000000001111111000000000;
			9'h0f5 : data = 24'b000000011111110000000000;
			9'h0f6 : data = 24'b000000111111100000000000;
			9'h0f7 : data = 24'b000001111111000000000000;
			9'h0f8 : data = 24'b000011111110000000000000;
			9'h0f9 : data = 24'b000111111100000000000000;
			9'h0fa : data = 24'b001111111000000000000000;
			9'h0fb : data = 24'b011111110000000000000000;
			9'h0fc : data = 24'b111111100000000000000000;
			9'h0fd : data = 24'b111111000000000000000000;
			9'h0fe : data = 24'b111110000000000000000000;
			9'h0ff : data = 24'b111100000000000000000000;
			
			// Eight
			9'h100 : data = 24'b000011111111111111110000;
			9'h101 : data = 24'b000111111111111111111000;
			9'h102 : data = 24'b001111111111111111111100;
			9'h103 : data = 24'b011111111111111111111110;
			9'h104 : data = 24'b111111100000000001111111;
			9'h105 : data = 24'b111111000000000000111111;
			9'h106 : data = 24'b111110000000000000011111;
			9'h107 : data = 24'b111100000000000000001111;
			9'h108 : data = 24'b111100000000000000001111;
			9'h109 : data = 24'b111100000000000000001111;
			9'h10a : data = 24'b111100000000000000001111;
			9'h10b : data = 24'b111110000000000000011111;
			9'h10c : data = 24'b111111000000000000111111;
			9'h10d : data = 24'b111111100000000001111111;
			9'h10e : data = 24'b011111111111111111111110;
			9'h10f : data = 24'b001111111111111111111100;
			9'h110 : data = 24'b000111111111111111111000;
			9'h111 : data = 24'b001111111111111111111100;
			9'h112 : data = 24'b011111100000000001111110;
			9'h113 : data = 24'b111111000000000000111111;
			9'h114 : data = 24'b111110000000000000011111;
			9'h115 : data = 24'b111100000000000000001111;
			9'h116 : data = 24'b111100000000000000001111;
			9'h117 : data = 24'b111100000000000000001111;
			9'h118 : data = 24'b111100000000000000001111;
			9'h119 : data = 24'b111110000000000000011111;
			9'h11a : data = 24'b111111000000000000111111;
			9'h11b : data = 24'b111111100000000001111111;
			9'h11c : data = 24'b011111111111111111111110;
			9'h11d : data = 24'b001111111111111111111100;
			9'h11e : data = 24'b000111111111111111111000;
			9'h11f : data = 24'b000011111111111111110000;
			
		endcase


endmodule
