`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    02:19:14 04/26/2012 
// Design Name: 
// Module Name:    turn_rom 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module turn_rom(
	 input wire clk,
	 input wire [5:0] addr,
	 output reg [79:0] data
    );
	 
	 // Registers used to access font ROM
	 reg [5:0] addr_reg;
	 reg [79:0] data_reg;
	 
	 always @ (posedge clk)
		addr_reg <= addr;
	 
	 // Font ROM
	 always @ *
		case (addr_reg)
			6'h00 : data = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
			6'h01 : data = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
			6'h02 : data = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
			6'h03 : data = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
			6'h04 : data = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
			6'h05 : data = 80'b00000000000100010000000000000000000000000000000000000000000000000000000000000000;
			6'h06 : data = 80'b00000010111100001110000000000000000000000000000000000000000000000000000000000000;
			6'h07 : data = 80'b00000001111111001110000000000000000000000000000000000000000000000000000000000000;
			6'h08 : data = 80'b00000001101110101100000000000000000000000000011000000000000000000000000000000000;
			6'h09 : data = 80'b00000000101111011000010111111000000001110011111101011101011000000000000000000000;
			6'h0a : data = 80'b00000000010111111000101111011110100111110011111000111111111000000000000000000000;
			6'h0b : data = 80'b00000000110111110000010110010111100101110010111000101111110000000000000000000000;
			6'h0c : data = 80'b00000000101011101000101110110111000101110110111001101110001000000000000000000000;
			6'h0d : data = 80'b00000000011111100000101110110111001101110111111001101110000000000000000000000000;
			6'h0e : data = 80'b00000000011111100000101110011111101111110111111000111110100000000000000000000000;
			6'h0f : data = 80'b00000000001111101000101110011111000111111011111000111110000000000000000000000000;
			6'h10 : data = 80'b00000000101111101000111110100111000111110111111000111111000000000000000000000000;
			6'h11 : data = 80'b00000000001111101000111111011110000111111111111000111111000000000000000000000000;
			6'h12 : data = 80'b00000000001111100000010111111000000111111001111000111111000000000000000000000000;
			6'h13 : data = 80'b00000000000000010000110000100010000000000000000100000001000000000000000000000000;
			6'h14 : data = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
			6'h15 : data = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
			6'h16 : data = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
			6'h17 : data = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
			6'h18 : data = 80'b00000000000000000000000000000010111000000000000000000000000000000000000000000000;
			6'h19 : data = 80'b00000000000000000000000111111111110000000000000000000000000000000000000000000000;
			6'h1a : data = 80'b00000000000000000000000111111111111000000000000000000000000000000000000000000000;
			6'h1b : data = 80'b00000000000000000000000100101110001000000000000100000000000000000000000000000000;
			6'h1c : data = 80'b00000000000000000000000001101110100000001000000001010011010110000110011101000000;
			6'h1d : data = 80'b00000000000000000000000010101110010001111100111101001111111110011110111110000000;
			6'h1e : data = 80'b00000000000000000000000010101110000001111110111100001011111100011111111111000000;
			6'h1f : data = 80'b00000000000000000000000000101110000001011100111100011011100100011111010111000000;
			6'h20 : data = 80'b00000000000000000000000000111110000011011100111100011111100100111110010111000000;
			6'h21 : data = 80'b00000000000000000000000000111110000011011101111100011111001000111111010111100000;
			6'h22 : data = 80'b00000000000000000000000000111110000001111100111110001111001000111111011111100000;
			6'h23 : data = 80'b00000000000000000000000000111110000001111100111110001111010000111111011111100000;
			6'h24 : data = 80'b00000000000000000000000000111110000001111111111110001111010000111110011111000000;
			6'h25 : data = 80'b00000000000000000000000000111110100000111110111110001111110000011110011110000000;
			6'h26 : data = 80'b00000000000000000000000001000000000001011101000001000000010000011100101000000000;
			6'h27 : data = 80'b00000000000000000000000001000000000000000000000000000000000000000000000000000000;
			6'h28 : data = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
			6'h29 : data = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
			6'h2a : data = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
			6'h2b : data = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
		endcase

endmodule
