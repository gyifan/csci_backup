`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Bucknell University
// Engineer: Yifan Ge, Alex Thompson
// 
// Create Date:    23:07:21 04/25/2012 
// Design Name: Memory Game Card Image
// Module Name:    card_rom 
// Project Name: Project 3 ELEC 340
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module card_rom(
	 input wire clk,
	 input wire [6:0] addr,
	 output reg [239:0] data
    );
	 
	 // Registers used to access font ROM
	 reg [6:0] addr_reg;
	 reg [239:0] data_reg;
	 
	 always @ (posedge clk)
		addr_reg <= addr;
	 
	 // Font ROM
	 always @ *
		case (addr_reg)
			// Thompson's face
			7'h00 : data = 240'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111011011011011011011011111111111111011111;
			7'h01 : data = 240'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111011011011011011011011111111111111011111;
			7'h02 : data = 240'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011011011011011011011011111111011111;
			7'h03 : data = 240'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011011011011011011011011111111011111;
			7'h04 : data = 240'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011011000000000000000000000000000000011111111111111111011111111111111111111111111111111111111111111011011011011011011011011011011111111111111011111;
			7'h05 : data = 240'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111011000000000000000000000000000000000000000000001011111011111011111111111111111111111111111111111111111111011011011011011011011011011011111111111011111;
			7'h06 : data = 240'b111111111111111111111111111111111111111111111111111111111111111111111111111111111011000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111011111011011011011011011011111111111111;
			7'h07 : data = 240'b111111111111111111111111111111111111111111111111111111111111111111111111111011001000000000000000000000000000000000000000000000000000000000000000000000011111111111111011111111111111111111111111111111111011111011011011011011011011111111111111;
			7'h08 : data = 240'b111111111111111111111111111111111111111111111111111111111111111111111111001000000000000000000000000000000000000000000000000000000000000000000000000000000111111111011111111111111111111111111111111111111111111011011011011011011011111111111111;
			7'h09 : data = 240'b111111111111111111111111111111111111111111111111111111111111111111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111011011011011011111011111111111111111111111011011011011111011011011011011111111;
			7'h0a : data = 240'b111111111111111111111111111111111111111111111111111111111111111001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111011011011011011011011011011111111111111011011011011011011011011011011111111;
			7'h0b : data = 240'b111111111111111111111111111111111111111111111111111111111111001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111011011011011011011111011011011011011011011011011011011111111011111111;
			7'h0c : data = 240'b111111111111111111111111111111111111111111111111111111111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011111111;
			7'h0d : data = 240'b111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111011011011011011011011011011011011011011011011011011011011011011111;
			7'h0e : data = 240'b111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111011011011011011011011011011011011011011011011011011111011111111;
			7'h0f : data = 240'b111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111011011011011011011011011011011011011011011011011011111111111111;
			7'h10 : data = 240'b111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011111111011111;
			7'h11 : data = 240'b111111111111111111111111111111111111111111111111011000000000000000000000000000000000000000000000100000000000000100100100110100000100000000000000000000000000000000000000000000001111011011011011011011011011011011011011011011011011011011011111;
			7'h12 : data = 240'b111111111111111111111111111111111111111111111111000000000000000000000000000000000000100000000100110100000100100110111110110100100110100100100100000000000000000000000000000000000111111011011011011011011011011011011011011011011011011011011111;
			7'h13 : data = 240'b111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000100100100100110110110110110110110110110110100110110100100000000000000000000000000000000011111011011011011011011011011011011011011011011011011011011111;
			7'h14 : data = 240'b111111111111111111111111111111111111111111111111000000000000000000000000100000100100100110110110110110110110110110110110110110110100110110110110110000000000000000000000000000000000111011011011011011011011011011011011011011011011011011011111;
			7'h15 : data = 240'b111111111111111111111111111111111111111111111111000000000000000000000100100110110110110110110110110110110111111111111110110110110110110110110110100000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011111;
			7'h16 : data = 240'b111111111111111111111111111111111111111111111001000000000000000000000100110110110110110110110110111111111111111111110111111111111110110110110110110100000000000000000000000000000000001111011011011011011011011011011011011011011011011011011111;
			7'h17 : data = 240'b111111111111111111111111111111111111111111111001000000000000000000100110110110110110110110110110111111111111111111111111111111111110110110110110110110100100100100100000000000000000000011011011011011011011011011011011011011011011011011011111;
			7'h18 : data = 240'b111111111111111111111111111111111111111111111001000000000000000000100100110110110110110110110110111111111111111111111111111111111111110110110110110110110110100100100100000000000000000011011011011011011011011011011011011011011011011011011111;
			7'h19 : data = 240'b111111111111111111111111111111111111111111111001000000000000000000100110110110110110110110110111111111111111110111111111111111111110110110110110110110110110110110100000000000000000000011011011011011011011011011011011011011011011011011011111;
			7'h1a : data = 240'b111111111111111111111111111111111111111111111011000000000000000000100110110110110110110110110110111110110111111111111111111111111111110110110110110110110110110110100100000000000000000011011011011011011011011011011011011011011011011011011111;
			7'h1b : data = 240'b111111111111111111111111111111111111111111111011000000000000000000100110110110110110110110110110110110111110110110111111111111111111110110110110110110110110110110100100000000000000000011011011011011011011011011011011011011011011011011011111;
			7'h1c : data = 240'b111111111111111111111111111111111111111111111011000000000000000000100110110110110110110110110111110111111111111111111111111111111111110110110110110110110110110110110100000000000000000011011011011011011011011011011011011011011011011011011111;
			7'h1d : data = 240'b111111111111111111111111111111111111111111111011000000000000000000110110110110110110110111111111111111111111111111111111111111111111110110110110110110110110110110100100000000000000000011011011011011011011011011011011011011011011011011011111;
			7'h1e : data = 240'b011111111111111111111111111111111111111111111011000000000000000100110110110110110110110111111111111111111111111111111111111111111111111111111110110110110110110110100100000000000000000011011011011011011011011011011011011011011011011011011111;
			7'h1f : data = 240'b011011111111111111111111111111111111111111111111000000000000000100110110110110110110110111111111111111111111111111111111111111111111111111111111111110110110110110110100000000000000000011011011011011011011011011011011011011011011011011011111;
			7'h20 : data = 240'b111111111111111111011111111111111111111111111111000000000000000100110110110110110110111111111111111111111111111111111111111111111111111111111111111111111111110110100100000000000000000011011011011011011011011011011011011011011011011011011111;
			7'h21 : data = 240'b111111111111111111111011111111011111111111111111000000000000000100110110110110110110110110110110110110110110110110111111111111111111111111111110110110110110110100110100000000000000000011011011011011011011011011011011011011011011011011011111;
			7'h22 : data = 240'b011011011011011011011011111111111111111111111101000000000000000100110110110111110110110110110100100100100100100110111111111111111111111110100100000000000000100100100100000000000000001011011011011011011011011011011011011011011011011011011111;
			7'h23 : data = 240'b011011011011011011011111111111111111111111100111111000000000100110110110110110110111111111111111111110100110110110110111111111111110110100100100100111111111111110100000000000000000000011011011011011011011011011011011011011011011011011011111;
			7'h24 : data = 240'b011011011011011011111111111111011111111111111100111000000000100110110110110111111111111110110100000100100100100100110110111111110110100000100100100000110110111111110100000000000000000001011011011011011011011011011011011011011011011011011111;
			7'h25 : data = 240'b011011011011011011111111111111011111111111111110111100000000110110110110111111111110100000000000000000100100110110100110111111110100000110100100000000000000000100110100100100000000000111111011011011011011011011011011011011011011011011011111;
			7'h26 : data = 240'b011011011011011111111111111011011111111111110110111110000000110110110111111111110100000100100000000111111110110111110110110111110100100110110111000000000110000000100100110100000000101111111011011011011011011011011011011011011011011011011111;
			7'h27 : data = 240'b111011011011011111111111011011011111111111110111110100000000110110111111111111110110110111111111110110110110111111110110110110110100100110111110111110100100100000100100111110000000111111111011011011011011011011011011011011011011011011011111;
			7'h28 : data = 240'b011011011011111111111111011011011111111111111111111111000000110110110111111111111111111111111111111110110110110110110110110110111110100100110110110110110110110110110110110110100000100111111011011011011011011011011011011011011011011011011111;
			7'h29 : data = 240'b011011011111111111111111011011011111111111111111111111000000110110110111111111111111111111111111111110110110110110110110110111111110100100110110110110110110110110111110110110100000100111011011011011011011011011011011011011011011011011011111;
			7'h2a : data = 240'b011011011011011011111011011011011111111111111100111111000000110110110111111111111111111111111111111111111111110110110110110110111110100100110110110110110110110110110110110100100000111111011011011011011011011011011011011011011011011011011111;
			7'h2b : data = 240'b011011011011011011011011011011011111111111110100110111100100100110110110111111111111111111111111111111111110110110110110110111110110100100100110110110110110110110110110110100100000111000011011011011011011011011011011011011011011011011011111;
			7'h2c : data = 240'b011011011011011011011111111011011111111111110110110111100100100110110111111111111111111111111111111111111110110110110110110111110110100100100110110110110110110110110110110100000000100000011011011011011011011011011011011011011011011011011111;
			7'h2d : data = 240'b011011111011011011011111111011011111111111110111111110100100100100110111111111111111111111111111111111111110110110110110110111111110100100100110110110110110110110110110110100000100000000011011011011011011011011011011011011011011011011011111;
			7'h2e : data = 240'b011011111111011011011111111111011111011100111111111111100100100100110110111111111111111111111111111111111111110110110110111111111111100100100110111111111111111110110110100100000110000000011011011011011011011011011011011011011011011011011111;
			7'h2f : data = 240'b011011011011011011011011111111011111011000111111111111100100100100110111111111111111111111111111111111111110100110110110111111111111110100100100111111111111111111110110100100000100000001011011011011011011011011011011011011011011011011011111;
			7'h30 : data = 240'b011011011011011011011011111011111111011000111111111111110000100100110110111111111111111111111111111111110110100110110110111111111111111100100100110111111111111111110110100100000100000001011011011011011011011011011011011011011011011011011111;
			7'h31 : data = 240'b011011011011011011011011011111111111011000000111111111110000100100110110111111110111111111111111111110110110110110110110111111111111111100100000110110110111111111111110100100000111000001011011011011011011011011011011011011011011011011011111;
			7'h32 : data = 240'b011011011011011011011011011011011111011000000000110110000100100100110110111110110111111111111111110110111111100110100100110110100110100000100100110110110111111111110110100000000111000001011011011011011011011011011011011011011011011011011111;
			7'h33 : data = 240'b011011111011011011011011011011011011011001000000000000000000000100100110111110110111111111111110110111111111111110110110100100100000000100100110110110110110110110110100100000000000000001011011011011011011011011011011011011011011011011011111;
			7'h34 : data = 240'b111111111111011011011011011011011011011001000000000000000000100100110110110111110110111111110110110111111111111111111111111110110111110100110100110110110110110110110100100000000000000011011011011011011011011011011011011011011011011011011111;
			7'h35 : data = 240'b011011111011011011011011011011011011011011000000000000000000100100100110110110110110110111110110111110111111111111111111111111111111110110100110110110110100110110110100100000000000000001011011011011011011011011011011011011011011011011011111;
			7'h36 : data = 240'b011011011011011011011011011011011011011011001000000000000000000100100110110110110110111110110110110110110110110111111111111111111111111110110100100110100100111110110100100000000000000001011011011011011011011011011011011011011011011011011111;
			7'h37 : data = 240'b011011011011011011011011011011011011011011011001000000000000000100110110110110110110111110110110110110110110110111111111111111111111110100100100000100110110111110110100100000000000000011011011011011011011011011011011011011011011011011011111;
			7'h38 : data = 240'b011011011011011011011011011011011011011011011011011011011000000000100110110110110110110110110110110000100100110100110100100100100100100100000000000111110110111110110100100000000000001011011011011011011011011011011011011011011011011011011111;
			7'h39 : data = 240'b011011011011011011011011111011011011011011011011111011011000000000100110110110110110110111110111111111100110110111111111111111111111100100100100110110110111111110110100000000001011011011011011011011011011011011011011011011011011011011011111;
			7'h3a : data = 240'b011011011011011011011011111011011011011011011011011011011001000000000100110110110110110111111111111111110100100100100100100100100100100100100100110110110111111110100100000000011011011011011011011011011011011011011011011011011011011011011111;
			7'h3b : data = 240'b011011111011011011011011111011011011011011011011011011011001000000000100110110110110110111110111111110110110110110110111111111111111100100100100100110110111110100100000000000011011011011011011011011011011011011011011011011011011011011011111;
			7'h3c : data = 240'b011011111011011011011011111011011011011011011011011111011011000000000000100110110110110110110110110110110110110110111111110111110110100110100100110110110111110100100000000000011011011011011011011011011011011011011011011011011011011011011111;
			7'h3d : data = 240'b011011011011011011011011111011011011011011011011011011111011000000000000100110110110110110111110110110110110110110111111111110110110110110100100110110110110100100000000000001011011011011011011011011011011011011011011011011011011011011011111;
			7'h3e : data = 240'b011011011011011011011011111011011011011011011011011011111111001000000000000100110110110110110110110110110110110110111110110110110110110110110110110110110110100000000000000001011011011011011011011011011011011011011011011011011011011011011111;
			7'h3f : data = 240'b011011011011011011011011011011011011011011011011011011011111011000000100000000100110110110110110110110110110110110110111111110110111110110110110110110110100000000000000000001011011011011011011011011011011011011011011011011011011011011011111;
			7'h40 : data = 240'b011011011011011011011011011011011011011011011011011011011111011000100100100000000110110110110110110110110110111110110111111110110110110110110110100100100000000000000000000001111011011011011011011011011011011011011011011011011011011011011111;
			7'h41 : data = 240'b011011011011011011011011011011011011011011011011011011011111111000100100100000000000110110110110111110110111110111111110110110110110110110110110100000000000000000000111111111011011011011011011011011011011011011011011011011011011011011011111;
			7'h42 : data = 240'b111011011011011011011011011011011111011011011011011011011111111000100110100100000000000100100100100110110110111111111111111111111110110110110100000000000000000000000111111000011011011011011011011011011011011011011011011011011011011011011111;
			7'h43 : data = 240'b111111011011011011011011111011011011011011011011011011111111111000100110110100100100000000100100100100110110110111111111111111111110110110100100000000000000000000000111111000000011011011011011011011011011011011011011011011011011011011011111;
			7'h44 : data = 240'b011011011011011011011011011011011011011011011011011011111111111000100100110110110100100000000000100100100110110110111111111111110110110110100000000000000000000000000111111111000011011011011011011011011011011011011011011011011011011011011111;
			7'h45 : data = 240'b011011011011011011011011011011011011011011011011011111111111001000100100110110110110110100000000000100000000100110110110110110110110100000000000000000000000000000000111001111000001111011011011011011011011011011011011011011011011011011011111;
			7'h46 : data = 240'b011011011011011011011011011011011011011011011011111111111001000000100100110110110110110110100100000000000000000000000000100000000000000000000000000000000000000000000111111000000000111011001011011011011011011011011011011011011011011011011111;
			7'h47 : data = 240'b011011011011011011011011011011011011011011011011111111111001000000100100110110110110110110110100110100000000000000000000000000000000000000000000000000000000000000000000111111111000111111001011011011011011011011011011011011011011011011011111;
			7'h48 : data = 240'b011011011011011011011011011011011011011011011011111111111001000111100100110110110110110110110110110110110110110100100100100000100100100100000000000000000000000000000000000000111000111111011011011011011011011011011011011011011011011011011111;
			7'h49 : data = 240'b011011011011011011011011011011011011011011011111111111111000111000100100100110110110110110110110110110110110110110110110110110110100100100000000000100100100000000000000000000111111111111011011011011011011011011011011011011011011011011011111;
			7'h4a : data = 240'b011011011011011011011011011011011011011011111111111111111111000000100100100110110110110110110110110110110110110110110111110111110110110100100000000100100100000000000000000000000111111111011111011011011011011011011011011011011011011011011111;
			7'h4b : data = 240'b011011011011011011011011011011011011011111111111111111111111000000000100100110110110110110110110110110110110110110110111111110110110110100100100100100100100000000000000000000000111111111111111111011111011011011011011011011011011011011011111;
			7'h4c : data = 240'b011011011011011011011011011011011011111111111111111111111111111000000100110110110110110110110110110110110110110110110110110110111100100100100100100100100100000000000000000000110111111111111111111111111111111011011011011011011011011011011111;
			7'h4d : data = 240'b011011011011011011011011011011111111111111111111111111111111111000000100110110110110110110110110110110110110110110110110110110110110100100100100100100100100100000000000000000111111111111111111111111111111111011111011011011011011011011011111;
			7'h4e : data = 240'b011011011011011011011011011011011111111111111111111111111111111111000100100110110110110110110110110110110110110110110110110110110100110100100110100100100100100000000000000100111111111111111111111111111111111111111111111111111011011011011111;
			7'h4f : data = 240'b011011011011011011011011011011011111111111111111111111111111111111111100110110110110110110110110110110110110110110111110110110110110110110110110110110110100100100000000000111111111111111111111111011111111111111111111111111111111111111011111;
		endcase

endmodule
